module sessions
