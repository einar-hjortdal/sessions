module sessions

// TODO test functions in jwt.v
fn test_init() {
	assert true
}
