module sessions